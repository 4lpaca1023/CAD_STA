//Generate the verilog at 2025-11-18T18:29:25 by iSTA.
module map9v3 (
N_0_,
N_1_,
N_2_,
N_3_,
N_4_,
N_5_,
N_6_,
N_7_,
N_8_,
clock,
counter_0_,
counter_1_,
counter_2_,
counter_3_,
counter_4_,
counter_5_,
counter_6_,
counter_7_,
done,
dp_0_,
dp_1_,
dp_2_,
dp_3_,
dp_4_,
dp_5_,
dp_6_,
dp_7_,
dp_8_,
reset,
sr_0_,
sr_1_,
sr_2_,
sr_3_,
sr_4_,
sr_5_,
sr_6_,
sr_7_,
start
);

input N_0_ ;
input N_1_ ;
input N_2_ ;
input N_3_ ;
input N_4_ ;
input N_5_ ;
input N_6_ ;
input N_7_ ;
input N_8_ ;
input clock ;
output counter_0_ ;
output counter_1_ ;
output counter_2_ ;
output counter_3_ ;
output counter_4_ ;
output counter_5_ ;
output counter_6_ ;
output counter_7_ ;
output done ;
output dp_0_ ;
output dp_1_ ;
output dp_2_ ;
output dp_3_ ;
output dp_4_ ;
output dp_5_ ;
output dp_6_ ;
output dp_7_ ;
output dp_8_ ;
input reset ;
output sr_0_ ;
output sr_1_ ;
output sr_2_ ;
output sr_3_ ;
output sr_4_ ;
output sr_5_ ;
output sr_6_ ;
output sr_7_ ;
input start ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire _136_ ;
wire _137_ ;
wire _138_ ;
wire _139_ ;
wire _140_ ;
wire _141_ ;
wire _142_ ;
wire _143_ ;
wire _144_ ;
wire _145_ ;
wire _146_ ;
wire _147_ ;
wire _148_ ;
wire _149_ ;
wire _150_ ;
wire _151_ ;
wire _152_ ;
wire _153_ ;
wire _154_ ;
wire _155_ ;
wire _156_ ;
wire _157_ ;
wire _158_ ;
wire _159_ ;
wire _160_ ;
wire _161_ ;
wire _162_ ;
wire _163_ ;
wire _164_ ;
wire _165_ ;
wire _166_ ;
wire startbuf ;
wire state_0_ ;
wire state_1_ ;
wire state_2_ ;
wire state_3_ ;
wire state_4_ ;
wire reset ;
wire start ;
wire N_4_ ;
wire N_5_ ;
wire N_0_ ;
wire N_1_ ;
wire N_2_ ;
wire N_3_ ;
wire N_6_ ;
wire N_7_ ;
wire N_8_ ;
wire counter_0_ ;
wire counter_1_ ;
wire counter_2_ ;
wire counter_3_ ;
wire counter_4_ ;
wire counter_5_ ;
wire counter_6_ ;
wire counter_7_ ;
wire done ;
wire dp_0_ ;
wire dp_1_ ;
wire dp_2_ ;
wire dp_3_ ;
wire dp_4_ ;
wire dp_5_ ;
wire dp_6_ ;
wire dp_7_ ;
wire dp_8_ ;
wire sr_0_ ;
wire sr_1_ ;
wire sr_2_ ;
wire sr_3_ ;
wire sr_4_ ;
wire sr_5_ ;
wire sr_6_ ;
wire sr_7_ ;
wire clock ;


INVX1 _167_ ( .A(reset ), .Y(_030_ ) );
INVX1 _168_ ( .A(state_3_ ), .Y(_031_ ) );
INVX1 _169_ ( .A(state_4_ ), .Y(_032_ ) );
INVX1 _170_ ( .A(state_1_ ), .Y(_033_ ) );
INVX1 _171_ ( .A(start ), .Y(_034_ ) );
INVX1 _172_ ( .A(state_0_ ), .Y(_035_ ) );
INVX1 _173_ ( .A(N_4_ ), .Y(_036_ ) );
INVX1 _174_ ( .A(N_5_ ), .Y(_037_ ) );
INVX1 _175_ ( .A(_149_ ), .Y(_038_ ) );
OR2X1 _176_ ( .A(_146_ ), .B(_145_ ), .Y(_039_ ) );
OR2X1 _177_ ( .A(_147_ ), .B(_039_ ), .Y(_040_ ) );
NOR2X1 _178_ ( .A(_144_ ), .B(_143_ ), .Y(_041_ ) );
NOR2X1 _179_ ( .A(_142_ ), .B(_141_ ), .Y(_042_ ) );
NAND2X1 _180_ ( .A(_041_ ), .B(_042_ ), .Y(_043_ ) );
OR2X1 _181_ ( .A(_040_ ), .B(_043_ ), .Y(_044_ ) );
OAI21X1 _182_ ( .A(_148_ ), .B(_044_ ), .C(state_3_ ), .Y(_045_ ) );
NAND2X1 _183_ ( .A(_035_ ), .B(_045_ ), .Y(_028_ ) );
NOR2X1 _184_ ( .A(startbuf ), .B(_034_ ), .Y(_046_ ) );
OAI21X1 _185_ ( .A(_033_ ), .B(_046_ ), .C(_032_ ), .Y(_029_ ) );
NAND3X1 _186_ ( .A(_031_ ), .B(state_2_ ), .C(_035_ ), .Y(_047_ ) );
MUX2X1 _187_ ( .A(_151_ ), .B(_159_ ), .S(_047_ ), .Y(_048_ ) );
INVX1 _188_ ( .A(_048_ ), .Y(_010_ ) );
MUX2X1 _189_ ( .A(_152_ ), .B(_160_ ), .S(_047_ ), .Y(_049_ ) );
INVX1 _190_ ( .A(_049_ ), .Y(_011_ ) );
MUX2X1 _191_ ( .A(_153_ ), .B(_161_ ), .S(_047_ ), .Y(_050_ ) );
INVX1 _192_ ( .A(_050_ ), .Y(_012_ ) );
MUX2X1 _193_ ( .A(_154_ ), .B(_162_ ), .S(_047_ ), .Y(_051_ ) );
INVX1 _194_ ( .A(_051_ ), .Y(_013_ ) );
MUX2X1 _195_ ( .A(_155_ ), .B(_163_ ), .S(_047_ ), .Y(_052_ ) );
INVX1 _196_ ( .A(_052_ ), .Y(_014_ ) );
MUX2X1 _197_ ( .A(_156_ ), .B(_164_ ), .S(_047_ ), .Y(_053_ ) );
INVX1 _198_ ( .A(_053_ ), .Y(_015_ ) );
MUX2X1 _199_ ( .A(_157_ ), .B(_165_ ), .S(_047_ ), .Y(_054_ ) );
INVX1 _200_ ( .A(_054_ ), .Y(_016_ ) );
MUX2X1 _201_ ( .A(_158_ ), .B(_166_ ), .S(_047_ ), .Y(_055_ ) );
INVX1 _202_ ( .A(_055_ ), .Y(_017_ ) );
MUX2X1 _203_ ( .A(_150_ ), .B(N_0_ ), .S(_047_ ), .Y(_056_ ) );
INVX1 _204_ ( .A(_056_ ), .Y(_009_ ) );
XOR2X1 _205_ ( .A(_164_ ), .B(_166_ ), .Y(_057_ ) );
XNOR2X1 _206_ ( .A(_162_ ), .B(_163_ ), .Y(_058_ ) );
XNOR2X1 _207_ ( .A(_057_ ), .B(_058_ ), .Y(_059_ ) );
OAI21X1 _208_ ( .A(state_3_ ), .B(_159_ ), .C(_035_ ), .Y(_060_ ) );
AOI21X1 _209_ ( .A(state_3_ ), .B(_059_ ), .C(_060_ ), .Y(_018_ ) );
NOR2X1 _210_ ( .A(state_3_ ), .B(_161_ ), .Y(_061_ ) );
OAI21X1 _211_ ( .A(_031_ ), .B(_160_ ), .C(_035_ ), .Y(_062_ ) );
NOR2X1 _212_ ( .A(_061_ ), .B(_062_ ), .Y(_020_ ) );
NOR2X1 _213_ ( .A(state_3_ ), .B(_162_ ), .Y(_063_ ) );
OAI21X1 _214_ ( .A(_031_ ), .B(_161_ ), .C(_035_ ), .Y(_064_ ) );
NOR2X1 _215_ ( .A(_063_ ), .B(_064_ ), .Y(_021_ ) );
NOR2X1 _216_ ( .A(state_3_ ), .B(_163_ ), .Y(_065_ ) );
OAI21X1 _217_ ( .A(_031_ ), .B(_162_ ), .C(_035_ ), .Y(_066_ ) );
NOR2X1 _218_ ( .A(_065_ ), .B(_066_ ), .Y(_022_ ) );
NOR2X1 _219_ ( .A(state_3_ ), .B(_164_ ), .Y(_067_ ) );
OAI21X1 _220_ ( .A(_031_ ), .B(_163_ ), .C(_035_ ), .Y(_068_ ) );
NOR2X1 _221_ ( .A(_067_ ), .B(_068_ ), .Y(_023_ ) );
NOR2X1 _222_ ( .A(state_3_ ), .B(_165_ ), .Y(_069_ ) );
OAI21X1 _223_ ( .A(_031_ ), .B(_164_ ), .C(_035_ ), .Y(_071_ ) );
NOR2X1 _224_ ( .A(_069_ ), .B(_071_ ), .Y(_024_ ) );
NOR2X1 _225_ ( .A(state_3_ ), .B(_166_ ), .Y(_074_ ) );
OAI21X1 _226_ ( .A(_031_ ), .B(_165_ ), .C(_035_ ), .Y(_076_ ) );
NOR2X1 _227_ ( .A(_074_ ), .B(_076_ ), .Y(_025_ ) );
XNOR2X1 _228_ ( .A(state_3_ ), .B(_141_ ), .Y(_079_ ) );
NAND2X1 _229_ ( .A(state_0_ ), .B(N_1_ ), .Y(_081_ ) );
OAI21X1 _230_ ( .A(state_0_ ), .B(_079_ ), .C(_081_ ), .Y(_000_ ) );
XOR2X1 _231_ ( .A(N_1_ ), .B(N_2_ ), .Y(_084_ ) );
NAND2X1 _232_ ( .A(state_3_ ), .B(_042_ ), .Y(_086_ ) );
OAI21X1 _233_ ( .A(_031_ ), .B(_141_ ), .C(_142_ ), .Y(_088_ ) );
NAND2X1 _234_ ( .A(_086_ ), .B(_088_ ), .Y(_090_ ) );
NAND2X1 _235_ ( .A(_035_ ), .B(_090_ ), .Y(_092_ ) );
OAI21X1 _236_ ( .A(_035_ ), .B(_084_ ), .C(_092_ ), .Y(_001_ ) );
AOI21X1 _237_ ( .A(N_1_ ), .B(N_2_ ), .C(N_3_ ), .Y(_095_ ) );
INVX1 _238_ ( .A(_095_ ), .Y(_097_ ) );
NAND3X1 _239_ ( .A(N_1_ ), .B(N_2_ ), .C(N_3_ ), .Y(_099_ ) );
NAND3X1 _240_ ( .A(state_0_ ), .B(_097_ ), .C(_099_ ), .Y(_101_ ) );
XOR2X1 _241_ ( .A(_143_ ), .B(_086_ ), .Y(_103_ ) );
OAI21X1 _242_ ( .A(state_0_ ), .B(_103_ ), .C(_101_ ), .Y(_002_ ) );
XNOR2X1 _243_ ( .A(_036_ ), .B(_095_ ), .Y(_106_ ) );
NAND3X1 _244_ ( .A(state_3_ ), .B(_041_ ), .C(_042_ ), .Y(_108_ ) );
OAI21X1 _245_ ( .A(_143_ ), .B(_086_ ), .C(_144_ ), .Y(_110_ ) );
AND2X1 _246_ ( .A(_035_ ), .B(_108_ ), .Y(_112_ ) );
AOI22X1 _247_ ( .A(state_0_ ), .B(_106_ ), .C(_110_ ), .D(_112_ ), .Y(_003_ ) );
NAND3X1 _248_ ( .A(_036_ ), .B(_037_ ), .C(_095_ ), .Y(_115_ ) );
OAI21X1 _249_ ( .A(N_4_ ), .B(_097_ ), .C(N_5_ ), .Y(_117_ ) );
NAND3X1 _250_ ( .A(state_0_ ), .B(_115_ ), .C(_117_ ), .Y(_119_ ) );
NOR2X1 _251_ ( .A(_145_ ), .B(_108_ ), .Y(_121_ ) );
XOR2X1 _252_ ( .A(_145_ ), .B(_108_ ), .Y(_123_ ) );
OAI21X1 _253_ ( .A(state_0_ ), .B(_123_ ), .C(_119_ ), .Y(_004_ ) );
AOI21X1 _254_ ( .A(N_6_ ), .B(_115_ ), .C(_035_ ), .Y(_125_ ) );
OAI21X1 _255_ ( .A(N_6_ ), .B(_115_ ), .C(_125_ ), .Y(_126_ ) );
XNOR2X1 _256_ ( .A(_146_ ), .B(_121_ ), .Y(_127_ ) );
OAI21X1 _257_ ( .A(state_0_ ), .B(_127_ ), .C(_126_ ), .Y(_005_ ) );
NOR3X1 _258_ ( .A(N_6_ ), .B(N_7_ ), .C(_115_ ), .Y(_128_ ) );
OAI21X1 _259_ ( .A(N_6_ ), .B(_115_ ), .C(N_7_ ), .Y(_129_ ) );
NAND2X1 _260_ ( .A(state_0_ ), .B(_129_ ), .Y(_130_ ) );
OR2X1 _261_ ( .A(_040_ ), .B(_108_ ), .Y(_131_ ) );
OAI21X1 _262_ ( .A(_039_ ), .B(_108_ ), .C(_147_ ), .Y(_132_ ) );
AND2X1 _263_ ( .A(_131_ ), .B(_132_ ), .Y(_133_ ) );
OAI22X1 _264_ ( .A(_128_ ), .B(_130_ ), .C(_133_ ), .D(state_0_ ), .Y(_006_ ) );
XOR2X1 _265_ ( .A(N_8_ ), .B(_128_ ), .Y(_134_ ) );
NOR2X1 _266_ ( .A(_148_ ), .B(_131_ ), .Y(_027_ ) );
XOR2X1 _267_ ( .A(_148_ ), .B(_131_ ), .Y(_135_ ) );
MUX2X1 _268_ ( .A(_134_ ), .B(_135_ ), .S(state_0_ ), .Y(_007_ ) );
NAND2X1 _269_ ( .A(_031_ ), .B(state_4_ ), .Y(_136_ ) );
OAI21X1 _270_ ( .A(state_2_ ), .B(_136_ ), .C(_038_ ), .Y(_137_ ) );
AND2X1 _271_ ( .A(_035_ ), .B(_137_ ), .Y(_008_ ) );
NOR2X1 _272_ ( .A(state_3_ ), .B(_160_ ), .Y(_138_ ) );
OAI21X1 _273_ ( .A(_031_ ), .B(_159_ ), .C(_035_ ), .Y(_139_ ) );
NOR2X1 _274_ ( .A(_138_ ), .B(_139_ ), .Y(_019_ ) );
NAND2X1 _275_ ( .A(state_1_ ), .B(_046_ ), .Y(_140_ ) );
INVX1 _276_ ( .A(_140_ ), .Y(_026_ ) );
INVX1 _277_ ( .A(reset ), .Y(_070_ ) );
INVX1 _278_ ( .A(reset ), .Y(_072_ ) );
INVX1 _279_ ( .A(reset ), .Y(_073_ ) );
INVX1 _280_ ( .A(reset ), .Y(_075_ ) );
INVX1 _281_ ( .A(reset ), .Y(_077_ ) );
INVX1 _282_ ( .A(reset ), .Y(_078_ ) );
INVX1 _283_ ( .A(reset ), .Y(_080_ ) );
INVX1 _284_ ( .A(reset ), .Y(_082_ ) );
INVX1 _285_ ( .A(reset ), .Y(_083_ ) );
INVX1 _286_ ( .A(reset ), .Y(_085_ ) );
INVX1 _287_ ( .A(reset ), .Y(_087_ ) );
INVX1 _288_ ( .A(reset ), .Y(_089_ ) );
INVX1 _289_ ( .A(reset ), .Y(_091_ ) );
INVX1 _290_ ( .A(reset ), .Y(_093_ ) );
INVX1 _291_ ( .A(reset ), .Y(_094_ ) );
INVX1 _292_ ( .A(reset ), .Y(_096_ ) );
INVX1 _293_ ( .A(reset ), .Y(_098_ ) );
INVX1 _294_ ( .A(reset ), .Y(_100_ ) );
INVX1 _295_ ( .A(reset ), .Y(_102_ ) );
INVX1 _296_ ( .A(reset ), .Y(_104_ ) );
INVX1 _297_ ( .A(reset ), .Y(_105_ ) );
INVX1 _298_ ( .A(reset ), .Y(_107_ ) );
INVX1 _299_ ( .A(reset ), .Y(_109_ ) );
INVX1 _300_ ( .A(reset ), .Y(_111_ ) );
INVX1 _301_ ( .A(reset ), .Y(_113_ ) );
INVX1 _302_ ( .A(reset ), .Y(_114_ ) );
INVX1 _303_ ( .A(reset ), .Y(_116_ ) );
INVX1 _304_ ( .A(reset ), .Y(_118_ ) );
INVX1 _305_ ( .A(reset ), .Y(_120_ ) );
INVX1 _306_ ( .A(reset ), .Y(_122_ ) );
INVX1 _307_ ( .A(reset ), .Y(_124_ ) );
BUFX2 _308_ ( .A(_141_ ), .Y(counter_0_ ) );
BUFX2 _309_ ( .A(_142_ ), .Y(counter_1_ ) );
BUFX2 _310_ ( .A(_143_ ), .Y(counter_2_ ) );
BUFX2 _311_ ( .A(_144_ ), .Y(counter_3_ ) );
BUFX2 _312_ ( .A(_145_ ), .Y(counter_4_ ) );
BUFX2 _313_ ( .A(_146_ ), .Y(counter_5_ ) );
BUFX2 _314_ ( .A(_147_ ), .Y(counter_6_ ) );
BUFX2 _315_ ( .A(_148_ ), .Y(counter_7_ ) );
BUFX2 _316_ ( .A(_149_ ), .Y(done ) );
BUFX2 _317_ ( .A(_150_ ), .Y(dp_0_ ) );
BUFX2 _318_ ( .A(_151_ ), .Y(dp_1_ ) );
BUFX2 _319_ ( .A(_152_ ), .Y(dp_2_ ) );
BUFX2 _320_ ( .A(_153_ ), .Y(dp_3_ ) );
BUFX2 _321_ ( .A(_154_ ), .Y(dp_4_ ) );
BUFX2 _322_ ( .A(_155_ ), .Y(dp_5_ ) );
BUFX2 _323_ ( .A(_156_ ), .Y(dp_6_ ) );
BUFX2 _324_ ( .A(_157_ ), .Y(dp_7_ ) );
BUFX2 _325_ ( .A(_158_ ), .Y(dp_8_ ) );
BUFX2 _326_ ( .A(_159_ ), .Y(sr_0_ ) );
BUFX2 _327_ ( .A(_160_ ), .Y(sr_1_ ) );
BUFX2 _328_ ( .A(_161_ ), .Y(sr_2_ ) );
BUFX2 _329_ ( .A(_162_ ), .Y(sr_3_ ) );
BUFX2 _330_ ( .A(_163_ ), .Y(sr_4_ ) );
BUFX2 _331_ ( .A(_164_ ), .Y(sr_5_ ) );
BUFX2 _332_ ( .A(_165_ ), .Y(sr_6_ ) );
BUFX2 _333_ ( .A(_166_ ), .Y(sr_7_ ) );
DFFSR _334_ ( .CLK(clock ), .D(_026_ ), .Q(state_0_ ), .R(1'b0 ), .S(_070_ ) );
DFFSR _335_ ( .CLK(clock ), .D(_029_ ), .Q(state_1_ ), .R(_072_ ), .S(1'b0 ) );
DFFSR _336_ ( .CLK(clock ), .D(_027_ ), .Q(state_2_ ), .R(_073_ ), .S(1'b0 ) );
DFFSR _337_ ( .CLK(clock ), .D(_028_ ), .Q(state_3_ ), .R(_075_ ), .S(1'b0 ) );
DFFSR _338_ ( .CLK(clock ), .D(state_2_ ), .Q(state_4_ ), .R(_077_ ), .S(1'b0 ) );
DFFSR _339_ ( .CLK(clock ), .D(_009_ ), .Q(_150_ ), .R(_078_ ), .S(1'b0 ) );
DFFSR _340_ ( .CLK(clock ), .D(_010_ ), .Q(_151_ ), .R(_080_ ), .S(1'b0 ) );
DFFSR _341_ ( .CLK(clock ), .D(_011_ ), .Q(_152_ ), .R(_082_ ), .S(1'b0 ) );
DFFSR _342_ ( .CLK(clock ), .D(_012_ ), .Q(_153_ ), .R(_083_ ), .S(1'b0 ) );
DFFSR _343_ ( .CLK(clock ), .D(_013_ ), .Q(_154_ ), .R(_085_ ), .S(1'b0 ) );
DFFSR _344_ ( .CLK(clock ), .D(_014_ ), .Q(_155_ ), .R(_087_ ), .S(1'b0 ) );
DFFSR _345_ ( .CLK(clock ), .D(_015_ ), .Q(_156_ ), .R(_089_ ), .S(1'b0 ) );
DFFSR _346_ ( .CLK(clock ), .D(_016_ ), .Q(_157_ ), .R(_091_ ), .S(1'b0 ) );
DFFSR _347_ ( .CLK(clock ), .D(_017_ ), .Q(_158_ ), .R(_093_ ), .S(1'b0 ) );
DFFSR _348_ ( .CLK(clock ), .D(_008_ ), .Q(_149_ ), .R(_094_ ), .S(1'b0 ) );
DFFSR _349_ ( .CLK(clock ), .D(_000_ ), .Q(_141_ ), .R(_096_ ), .S(1'b0 ) );
DFFSR _350_ ( .CLK(clock ), .D(_001_ ), .Q(_142_ ), .R(_098_ ), .S(1'b0 ) );
DFFSR _351_ ( .CLK(clock ), .D(_002_ ), .Q(_143_ ), .R(_100_ ), .S(1'b0 ) );
DFFSR _352_ ( .CLK(clock ), .D(_003_ ), .Q(_144_ ), .R(_102_ ), .S(1'b0 ) );
DFFSR _353_ ( .CLK(clock ), .D(_004_ ), .Q(_145_ ), .R(_104_ ), .S(1'b0 ) );
DFFSR _354_ ( .CLK(clock ), .D(_005_ ), .Q(_146_ ), .R(_105_ ), .S(1'b0 ) );
DFFSR _355_ ( .CLK(clock ), .D(_006_ ), .Q(_147_ ), .R(_107_ ), .S(1'b0 ) );
DFFSR _356_ ( .CLK(clock ), .D(_007_ ), .Q(_148_ ), .R(_109_ ), .S(1'b0 ) );
DFFSR _357_ ( .CLK(clock ), .D(_018_ ), .Q(_159_ ), .R(_111_ ), .S(1'b0 ) );
DFFSR _358_ ( .CLK(clock ), .D(_019_ ), .Q(_160_ ), .R(_113_ ), .S(1'b0 ) );
DFFSR _359_ ( .CLK(clock ), .D(_020_ ), .Q(_161_ ), .R(_114_ ), .S(1'b0 ) );
DFFSR _360_ ( .CLK(clock ), .D(_021_ ), .Q(_162_ ), .R(_116_ ), .S(1'b0 ) );
DFFSR _361_ ( .CLK(clock ), .D(_022_ ), .Q(_163_ ), .R(_118_ ), .S(1'b0 ) );
DFFSR _362_ ( .CLK(clock ), .D(_023_ ), .Q(_164_ ), .R(_120_ ), .S(1'b0 ) );
DFFSR _363_ ( .CLK(clock ), .D(_024_ ), .Q(_165_ ), .R(_122_ ), .S(1'b0 ) );
DFFSR _364_ ( .CLK(clock ), .D(_025_ ), .Q(_166_ ), .R(_124_ ), .S(1'b0 ) );
DFFSR _365_ ( .CLK(clock ), .D(start ), .Q(startbuf ), .R(_030_ ), .S(1'b0 ) );

endmodule
